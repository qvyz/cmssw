
--- Algo template Generated from gt-algorithm: p2gt_algos.vhdl
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.all;

use work.ipbus.all;
use work.emp_data_types.all;
use work.emp_project_decl.all;

use work.emp_device_decl.all;
use work.emp_ttc_decl.all;

use work.common_pkg.all;

entity p2gt_algos is
  generic (
    cut_offset                                 : natural := 0
  );
  port (
    clk                                        : in std_logic; -- ipbus signals
    rst                                        : in std_logic;
    ipb_in                                     : in ipb_wbus;
    ipb_out                                    : out ipb_rbus;
    clk_algo                                   : in std_logic;
    rst_algo                                   : in std_logic;
    clk40                                      : in std_logic;
    rst40                                      : in std_logic;
    objects_valid                              : in std_logic;
    objects                                    : in t_obj_array(NUM_OBJ_TYPES-1 downto 0);
    algo_bits_valid_out                        : out std_logic;
    algo_bits_out                              : out std_logic_vector(NUM_ALGOS_IN_SRL-1 downto 0)
  );

end p2gt_algos;

architecture rtl of p2gt_algos is
  signal algo_bits_int, algo_bits_int2         : std_logic_vector(NUM_ALGOS_IN_SRL-1 downto 0);
  signal algo_bits_srl1_int                    : std_logic_vector(NUM_ALGOS_IN_SRL-1 downto 0);
  signal algo_bits_srl2_int                    : std_logic_vector(NUM_ALGOS_IN_SRL-1 downto 0);

  signal delayed_valid_to_payload : std_logic_vector(ALGO_REPLICATION_IN_SRL-1 downto 0);
  signal delayed_valid_buffer     : std_logic_vector(ALGO_LATENCY-1 downto 0);  -- TODO: 1 tick used for registering algo bits.
signal HLT_path0 : std_logic;
signal HLT_path1 : std_logic;
signal HLT_path2 : std_logic;
signal HLT_path3 : std_logic;
signal HLT_path4 : std_logic;
signal HLT_path5 : std_logic;
signal HLT_path6 : std_logic;
signal HLT_path7 : std_logic;
signal HLT_path8 : std_logic;
signal HLT_path9 : std_logic;
signal HLT_path10 : std_logic;
signal HLT_path11 : std_logic;
signal HLT_path12 : std_logic;
signal HLT_path13 : std_logic;
signal HLT_path14 : std_logic;
signal HLT_path15 : std_logic;
signal HLT_path16 : std_logic;
signal HLT_path17 : std_logic;
signal HLT_path18 : std_logic;
signal HLT_path19 : std_logic;
signal test_trf : std_logic;
signal test_trf1 : std_logic;
signal test_trf2 : std_logic;
signal test_trf3 : std_logic;




begin
  ipb_out <= IPB_RBUS_NULL;

  delayed_valid_buffer(0) <= delayed_valid_to_payload(0);

  process(clk_algo)
  begin
    if rising_edge(clk_algo) then
      delayed_valid_buffer(delayed_valid_buffer'high downto 1) <= delayed_valid_buffer(delayed_valid_buffer'high-1 downto 0);
    end if;
  end process;





  algos : for i in 0 to ALGO_REPLICATION_IN_SRL-1 generate
    signal delayed_objects_tmp : t_delayed_obj_array(0 to 4);
    signal delayed_objects     : t_delayed_obj_array(0 to 4);
    signal delayed_valid_tmp   : std_logic_vector(0 to 4);
    signal delayed_valid       : std_logic_vector(0 to 4);

    ATTRIBUTE max_fanout                    : integer;
    ATTRIBUTE max_fanout of delayed_objects : signal is 10;
    ATTRIBUTE max_fanout of delayed_valid   : signal is 10;
  begin 
    object_delay : entity work.p2gt_objectDelay
    port map (
      clk_algo        => clk_algo,
      rst_algo        => rst_algo,
      objects_valid   => objects_valid,
      objects         => objects,
      delayed_objects => delayed_objects_tmp,
      delayed_valid   => delayed_valid_tmp
    );



    reg_objects : process(clk_algo)
    begin
      if rising_edge(clk_algo) then
        delayed_objects <= delayed_objects_tmp;
        delayed_valid   <= delayed_valid_tmp;
      end if;
    end process reg_objects;

  delayed_valid_to_payload(i) <= delayed_valid(BX_ZERO);



HLTtestfilt0 : entity work.p2gt_doubleObjCond
generic map (
different_objects => true,
pT1_cut=> to_unsigned(5,14),
pT2_cut=> to_unsigned(7,14),
minEta1_cut=> to_signed(3,12),
minEta2_cut=> to_signed(3,12),
maxEta1_cut=> to_signed(36,12),
maxEta2_cut=> to_signed(50,12),
ss_cut => true 
)

port map (
clk           => clk, -- ipbus signals
rst           => rst,
ipb_in        => ipb_in,
ipb_out       => open,
clk_algo => clk_algo,
rst_algo => rst_algo,
objects_valid => delayed_valid(BX_ZERO),
object1=>delayed_objects(BX_ZERO)(MU_SLOT),
object2=>delayed_objects(BX_ZERO)(ELECTRON_SLOT),
algo_bit_out =>HLT_path0
      );




HLTtestfilt1 : entity work.p2gt_doubleObjCond
generic map (
different_objects => true,
pT1_cut=> to_unsigned(6,14),
pT2_cut=> to_unsigned(7,14),
minEta1_cut=> to_signed(3,12),
minEta2_cut=> to_signed(3,12),
maxEta1_cut=> to_signed(36,12),
maxEta2_cut=> to_signed(50,12),
ss_cut => true 
)

port map (
clk           => clk, -- ipbus signals
rst           => rst,
ipb_in        => ipb_in,
ipb_out       => open,
clk_algo => clk_algo,
rst_algo => rst_algo,
objects_valid => delayed_valid(BX_ZERO),
object1=>delayed_objects(BX_ZERO)(MU_SLOT),
object2=>delayed_objects(BX_ZERO)(ELECTRON_SLOT),
algo_bit_out =>HLT_path1
      );




HLTtestfilt2 : entity work.p2gt_doubleObjCond
generic map (
different_objects => true,
pT1_cut=> to_unsigned(7,14),
pT2_cut=> to_unsigned(7,14),
minEta1_cut=> to_signed(3,12),
minEta2_cut=> to_signed(3,12),
maxEta1_cut=> to_signed(36,12),
maxEta2_cut=> to_signed(50,12),
ss_cut => true 
)

port map (
clk           => clk, -- ipbus signals
rst           => rst,
ipb_in        => ipb_in,
ipb_out       => open,
clk_algo => clk_algo,
rst_algo => rst_algo,
objects_valid => delayed_valid(BX_ZERO),
object1=>delayed_objects(BX_ZERO)(MU_SLOT),
object2=>delayed_objects(BX_ZERO)(ELECTRON_SLOT),
algo_bit_out =>HLT_path2
      );




HLTtestfilt3 : entity work.p2gt_doubleObjCond
generic map (
different_objects => true,
pT1_cut=> to_unsigned(8,14),
pT2_cut=> to_unsigned(7,14),
minEta1_cut=> to_signed(3,12),
minEta2_cut=> to_signed(3,12),
maxEta1_cut=> to_signed(36,12),
maxEta2_cut=> to_signed(50,12),
ss_cut => true 
)

port map (
clk           => clk, -- ipbus signals
rst           => rst,
ipb_in        => ipb_in,
ipb_out       => open,
clk_algo => clk_algo,
rst_algo => rst_algo,
objects_valid => delayed_valid(BX_ZERO),
object1=>delayed_objects(BX_ZERO)(MU_SLOT),
object2=>delayed_objects(BX_ZERO)(ELECTRON_SLOT),
algo_bit_out =>HLT_path3
      );




HLTtestfilt4 : entity work.p2gt_doubleObjCond
generic map (
different_objects => true,
pT1_cut=> to_unsigned(9,14),
pT2_cut=> to_unsigned(7,14),
minEta1_cut=> to_signed(3,12),
minEta2_cut=> to_signed(3,12),
maxEta1_cut=> to_signed(36,12),
maxEta2_cut=> to_signed(50,12),
ss_cut => true 
)

port map (
clk           => clk, -- ipbus signals
rst           => rst,
ipb_in        => ipb_in,
ipb_out       => open,
clk_algo => clk_algo,
rst_algo => rst_algo,
objects_valid => delayed_valid(BX_ZERO),
object1=>delayed_objects(BX_ZERO)(MU_SLOT),
object2=>delayed_objects(BX_ZERO)(ELECTRON_SLOT),
algo_bit_out =>HLT_path4
      );




HLTtestfilt5 : entity work.p2gt_doubleObjCond
generic map (
different_objects => true,
pT1_cut=> to_unsigned(10,14),
pT2_cut=> to_unsigned(7,14),
minEta1_cut=> to_signed(3,12),
minEta2_cut=> to_signed(3,12),
maxEta1_cut=> to_signed(36,12),
maxEta2_cut=> to_signed(50,12),
ss_cut => true 
)

port map (
clk           => clk, -- ipbus signals
rst           => rst,
ipb_in        => ipb_in,
ipb_out       => open,
clk_algo => clk_algo,
rst_algo => rst_algo,
objects_valid => delayed_valid(BX_ZERO),
object1=>delayed_objects(BX_ZERO)(MU_SLOT),
object2=>delayed_objects(BX_ZERO)(ELECTRON_SLOT),
algo_bit_out =>HLT_path5
      );




HLTtestfilt6 : entity work.p2gt_doubleObjCond
generic map (
different_objects => true,
pT1_cut=> to_unsigned(11,14),
pT2_cut=> to_unsigned(7,14),
minEta1_cut=> to_signed(3,12),
minEta2_cut=> to_signed(3,12),
maxEta1_cut=> to_signed(36,12),
maxEta2_cut=> to_signed(50,12),
ss_cut => true 
)

port map (
clk           => clk, -- ipbus signals
rst           => rst,
ipb_in        => ipb_in,
ipb_out       => open,
clk_algo => clk_algo,
rst_algo => rst_algo,
objects_valid => delayed_valid(BX_ZERO),
object1=>delayed_objects(BX_ZERO)(MU_SLOT),
object2=>delayed_objects(BX_ZERO)(ELECTRON_SLOT),
algo_bit_out =>HLT_path6
      );




HLTtestfilt7 : entity work.p2gt_doubleObjCond
generic map (
different_objects => true,
pT1_cut=> to_unsigned(12,14),
pT2_cut=> to_unsigned(7,14),
minEta1_cut=> to_signed(3,12),
minEta2_cut=> to_signed(3,12),
maxEta1_cut=> to_signed(36,12),
maxEta2_cut=> to_signed(50,12),
ss_cut => true 
)

port map (
clk           => clk, -- ipbus signals
rst           => rst,
ipb_in        => ipb_in,
ipb_out       => open,
clk_algo => clk_algo,
rst_algo => rst_algo,
objects_valid => delayed_valid(BX_ZERO),
object1=>delayed_objects(BX_ZERO)(MU_SLOT),
object2=>delayed_objects(BX_ZERO)(ELECTRON_SLOT),
algo_bit_out =>HLT_path7
      );




HLTtestfilt8 : entity work.p2gt_doubleObjCond
generic map (
different_objects => true,
pT1_cut=> to_unsigned(13,14),
pT2_cut=> to_unsigned(7,14),
minEta1_cut=> to_signed(3,12),
minEta2_cut=> to_signed(3,12),
maxEta1_cut=> to_signed(36,12),
maxEta2_cut=> to_signed(50,12),
ss_cut => true 
)

port map (
clk           => clk, -- ipbus signals
rst           => rst,
ipb_in        => ipb_in,
ipb_out       => open,
clk_algo => clk_algo,
rst_algo => rst_algo,
objects_valid => delayed_valid(BX_ZERO),
object1=>delayed_objects(BX_ZERO)(MU_SLOT),
object2=>delayed_objects(BX_ZERO)(ELECTRON_SLOT),
algo_bit_out =>HLT_path8
      );




HLTtestfilt9 : entity work.p2gt_doubleObjCond
generic map (
different_objects => true,
pT1_cut=> to_unsigned(14,14),
pT2_cut=> to_unsigned(7,14),
minEta1_cut=> to_signed(3,12),
minEta2_cut=> to_signed(3,12),
maxEta1_cut=> to_signed(36,12),
maxEta2_cut=> to_signed(50,12),
ss_cut => true 
)

port map (
clk           => clk, -- ipbus signals
rst           => rst,
ipb_in        => ipb_in,
ipb_out       => open,
clk_algo => clk_algo,
rst_algo => rst_algo,
objects_valid => delayed_valid(BX_ZERO),
object1=>delayed_objects(BX_ZERO)(MU_SLOT),
object2=>delayed_objects(BX_ZERO)(ELECTRON_SLOT),
algo_bit_out =>HLT_path9
      );




HLTtestfilt10 : entity work.p2gt_doubleObjCond
generic map (
different_objects => true,
pT1_cut=> to_unsigned(15,14),
pT2_cut=> to_unsigned(7,14),
minEta1_cut=> to_signed(3,12),
minEta2_cut=> to_signed(3,12),
maxEta1_cut=> to_signed(36,12),
maxEta2_cut=> to_signed(50,12),
ss_cut => true 
)

port map (
clk           => clk, -- ipbus signals
rst           => rst,
ipb_in        => ipb_in,
ipb_out       => open,
clk_algo => clk_algo,
rst_algo => rst_algo,
objects_valid => delayed_valid(BX_ZERO),
object1=>delayed_objects(BX_ZERO)(MU_SLOT),
object2=>delayed_objects(BX_ZERO)(ELECTRON_SLOT),
algo_bit_out =>HLT_path10
      );




HLTtestfilt11 : entity work.p2gt_doubleObjCond
generic map (
different_objects => true,
pT1_cut=> to_unsigned(16,14),
pT2_cut=> to_unsigned(7,14),
minEta1_cut=> to_signed(3,12),
minEta2_cut=> to_signed(3,12),
maxEta1_cut=> to_signed(36,12),
maxEta2_cut=> to_signed(50,12),
ss_cut => true 
)

port map (
clk           => clk, -- ipbus signals
rst           => rst,
ipb_in        => ipb_in,
ipb_out       => open,
clk_algo => clk_algo,
rst_algo => rst_algo,
objects_valid => delayed_valid(BX_ZERO),
object1=>delayed_objects(BX_ZERO)(MU_SLOT),
object2=>delayed_objects(BX_ZERO)(ELECTRON_SLOT),
algo_bit_out =>HLT_path11
      );




HLTtestfilt12 : entity work.p2gt_doubleObjCond
generic map (
different_objects => true,
pT1_cut=> to_unsigned(17,14),
pT2_cut=> to_unsigned(7,14),
minEta1_cut=> to_signed(3,12),
minEta2_cut=> to_signed(3,12),
maxEta1_cut=> to_signed(36,12),
maxEta2_cut=> to_signed(50,12),
ss_cut => true 
)

port map (
clk           => clk, -- ipbus signals
rst           => rst,
ipb_in        => ipb_in,
ipb_out       => open,
clk_algo => clk_algo,
rst_algo => rst_algo,
objects_valid => delayed_valid(BX_ZERO),
object1=>delayed_objects(BX_ZERO)(MU_SLOT),
object2=>delayed_objects(BX_ZERO)(ELECTRON_SLOT),
algo_bit_out =>HLT_path12
      );




HLTtestfilt13 : entity work.p2gt_doubleObjCond
generic map (
different_objects => true,
pT1_cut=> to_unsigned(18,14),
pT2_cut=> to_unsigned(7,14),
minEta1_cut=> to_signed(3,12),
minEta2_cut=> to_signed(3,12),
maxEta1_cut=> to_signed(36,12),
maxEta2_cut=> to_signed(50,12),
ss_cut => true 
)

port map (
clk           => clk, -- ipbus signals
rst           => rst,
ipb_in        => ipb_in,
ipb_out       => open,
clk_algo => clk_algo,
rst_algo => rst_algo,
objects_valid => delayed_valid(BX_ZERO),
object1=>delayed_objects(BX_ZERO)(MU_SLOT),
object2=>delayed_objects(BX_ZERO)(ELECTRON_SLOT),
algo_bit_out =>HLT_path13
      );




HLTtestfilt14 : entity work.p2gt_doubleObjCond
generic map (
different_objects => true,
pT1_cut=> to_unsigned(19,14),
pT2_cut=> to_unsigned(7,14),
minEta1_cut=> to_signed(3,12),
minEta2_cut=> to_signed(3,12),
maxEta1_cut=> to_signed(36,12),
maxEta2_cut=> to_signed(50,12),
ss_cut => true 
)

port map (
clk           => clk, -- ipbus signals
rst           => rst,
ipb_in        => ipb_in,
ipb_out       => open,
clk_algo => clk_algo,
rst_algo => rst_algo,
objects_valid => delayed_valid(BX_ZERO),
object1=>delayed_objects(BX_ZERO)(MU_SLOT),
object2=>delayed_objects(BX_ZERO)(ELECTRON_SLOT),
algo_bit_out =>HLT_path14
      );




HLTtestfilt15 : entity work.p2gt_doubleObjCond
generic map (
different_objects => true,
pT1_cut=> to_unsigned(20,14),
pT2_cut=> to_unsigned(7,14),
minEta1_cut=> to_signed(3,12),
minEta2_cut=> to_signed(3,12),
maxEta1_cut=> to_signed(36,12),
maxEta2_cut=> to_signed(50,12),
ss_cut => true 
)

port map (
clk           => clk, -- ipbus signals
rst           => rst,
ipb_in        => ipb_in,
ipb_out       => open,
clk_algo => clk_algo,
rst_algo => rst_algo,
objects_valid => delayed_valid(BX_ZERO),
object1=>delayed_objects(BX_ZERO)(MU_SLOT),
object2=>delayed_objects(BX_ZERO)(ELECTRON_SLOT),
algo_bit_out =>HLT_path15
      );




HLTtestfilt16 : entity work.p2gt_doubleObjCond
generic map (
different_objects => true,
pT1_cut=> to_unsigned(21,14),
pT2_cut=> to_unsigned(7,14),
minEta1_cut=> to_signed(3,12),
minEta2_cut=> to_signed(3,12),
maxEta1_cut=> to_signed(36,12),
maxEta2_cut=> to_signed(50,12),
ss_cut => true 
)

port map (
clk           => clk, -- ipbus signals
rst           => rst,
ipb_in        => ipb_in,
ipb_out       => open,
clk_algo => clk_algo,
rst_algo => rst_algo,
objects_valid => delayed_valid(BX_ZERO),
object1=>delayed_objects(BX_ZERO)(MU_SLOT),
object2=>delayed_objects(BX_ZERO)(ELECTRON_SLOT),
algo_bit_out =>HLT_path16
      );




HLTtestfilt17 : entity work.p2gt_doubleObjCond
generic map (
different_objects => true,
pT1_cut=> to_unsigned(22,14),
pT2_cut=> to_unsigned(7,14),
minEta1_cut=> to_signed(3,12),
minEta2_cut=> to_signed(3,12),
maxEta1_cut=> to_signed(36,12),
maxEta2_cut=> to_signed(50,12),
ss_cut => true 
)

port map (
clk           => clk, -- ipbus signals
rst           => rst,
ipb_in        => ipb_in,
ipb_out       => open,
clk_algo => clk_algo,
rst_algo => rst_algo,
objects_valid => delayed_valid(BX_ZERO),
object1=>delayed_objects(BX_ZERO)(MU_SLOT),
object2=>delayed_objects(BX_ZERO)(ELECTRON_SLOT),
algo_bit_out =>HLT_path17
      );




HLTtestfilt18 : entity work.p2gt_doubleObjCond
generic map (
different_objects => true,
pT1_cut=> to_unsigned(23,14),
pT2_cut=> to_unsigned(7,14),
minEta1_cut=> to_signed(3,12),
minEta2_cut=> to_signed(3,12),
maxEta1_cut=> to_signed(36,12),
maxEta2_cut=> to_signed(50,12),
ss_cut => true 
)

port map (
clk           => clk, -- ipbus signals
rst           => rst,
ipb_in        => ipb_in,
ipb_out       => open,
clk_algo => clk_algo,
rst_algo => rst_algo,
objects_valid => delayed_valid(BX_ZERO),
object1=>delayed_objects(BX_ZERO)(MU_SLOT),
object2=>delayed_objects(BX_ZERO)(ELECTRON_SLOT),
algo_bit_out =>HLT_path18
      );




HLTtestfilt19 : entity work.p2gt_doubleObjCond
generic map (
different_objects => true,
pT1_cut=> to_unsigned(24,14),
pT2_cut=> to_unsigned(7,14),
minEta1_cut=> to_signed(3,12),
minEta2_cut=> to_signed(3,12),
maxEta1_cut=> to_signed(36,12),
maxEta2_cut=> to_signed(50,12),
ss_cut => true 
)

port map (
clk           => clk, -- ipbus signals
rst           => rst,
ipb_in        => ipb_in,
ipb_out       => open,
clk_algo => clk_algo,
rst_algo => rst_algo,
objects_valid => delayed_valid(BX_ZERO),
object1=>delayed_objects(BX_ZERO)(MU_SLOT),
object2=>delayed_objects(BX_ZERO)(ELECTRON_SLOT),
algo_bit_out =>HLT_path19
      );





  end generate;

  reg_outputs : process(clk_algo)  -- Register on algo clk for one BX
  begin
    if rising_edge(clk_algo) then 
	algo_bits_int2(0) <= HLT_path0 ;
	algo_bits_int2(1) <= HLT_path1 ;
	algo_bits_int2(2) <= HLT_path2 ;
	algo_bits_int2(3) <= HLT_path3 ;
	algo_bits_int2(4) <= HLT_path4 ;
	algo_bits_int2(5) <= HLT_path5 ;
	algo_bits_int2(6) <= HLT_path6 ;
	algo_bits_int2(7) <= HLT_path7 ;
	algo_bits_int2(8) <= HLT_path8 ;
	algo_bits_int2(9) <= HLT_path9 ;
	algo_bits_int2(10) <= HLT_path10 ;
	algo_bits_int2(11) <= HLT_path11 ;
	algo_bits_int2(12) <= HLT_path12 ;
	algo_bits_int2(13) <= HLT_path13 ;
	algo_bits_int2(14) <= HLT_path14 ;
	algo_bits_int2(15) <= HLT_path15 ;
	algo_bits_int2(16) <= HLT_path16 ;
	algo_bits_int2(17) <= HLT_path17 ;
	algo_bits_int2(18) <= HLT_path18 ;
	algo_bits_int2(19) <= HLT_path19 ;
	algo_bits_int2(20) <= HLT_path0 OR HLT_path19 ;
	algo_bits_int2(21) <= HLT_path1 OR HLT_path18 ;
	algo_bits_int2(22) <= HLT_path2 OR HLT_path17 ;
	algo_bits_int2(23) <= HLT_path3 OR HLT_path16 ;

        algo_bits_out <= algo_bits_int2;
    end if;
  end process;
  algo_bits_valid_out <= delayed_valid_buffer(delayed_valid_buffer'high);

end rtl;
